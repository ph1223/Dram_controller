task send_inputs();

endtask

task update_score_board();

endtask

task run_agent();

endtask