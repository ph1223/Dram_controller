`include "define.sv"

import user_types::*;
class ScoreBoard();
    data_t



endclass